module Q1_a(A, B, C, D, f);
input A, B, C, D;
output f;
assign f = (A&D)|C;
endmodule
